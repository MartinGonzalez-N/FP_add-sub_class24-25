package global_params;
    parameter int MANT_BITS = 23;
    parameter int EXP_BITS   = 8;  // Bits del exponente
    parameter int BIAS       = 127; // Sesgo del exponente para formato simple
endpackage
