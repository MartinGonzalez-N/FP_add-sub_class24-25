`define MID_VAl 32'h3f800000
`define INF 32'h7f800000
`define NEG_INF 32'hff800000
`define NAN 32'h7fc00000
`define MAX_POS 32'h7f7fffff
`define MIN_POS 32'h00800000 //Normalized
`define MIN_POS_DENORM 32'h00000001 //Denormalized
`define MAX_NEG 32'hff7fffff
`define MIN_NEG 32'h80800000 //Normalized
`define MIN_NEG_DENORM 32'h80000001 //Denormalized
`define CICLES 1000
`define WIDTH 32
`define ADD_SEL 1
`define SUB_SEL 0
`define SIGN_MASK 32'h80000000
`define EXP_MASK 32'h7f800000
`define MANT_MASK 32'h007fffff
`define NEG_INF 32'hff800000
`define ZERO 32'h00000000
`define ZERO_BIT 1'b0 
`define ONE_BIT 1'b1

